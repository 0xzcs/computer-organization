LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY ALU IS
PORT(
	A:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	B:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	S1,S0:IN STD_LOGIC;
	BCDOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	CF,ZF:OUT STD_LOGIC
	);
END ALU;
ARCHITECTURE A OF ALU IS
SIGNAL AA,BB,TEMP:STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
	PROCESS
	BEGIN
		IF(S1='0' AND S0='1') THEN
			BCDOUT <=A-B;
			IF(A<B) THEN
				CF<='1';
				ZF<='0';
			ELSIF(A=B) THEN
				CF<='0';
				ZF<='1';
			ELSE
				CF<='0';
				ZF<='0';
			END IF;
		ELSIF(S1='1' AND S0='0') THEN
			AA<='0'&A;
			BB<='0'&B;
			TEMP<=AA+BB;
			BCDOUT<=TEMP(7 DOWNTO 0);
			CF<=TEMP(8);
			IF(TEMP="100000000" OR TEMP ="000000000") THEN
				ZF<='1';
			ELSE
				ZF<='0';
			END IF;
		ELSIF(S1='1' AND S0='1') THEN
			BCDOUT<='0'&A(7 DOWNTO 1);
			CF<=A(0);
		ELSE 
			BCDOUT<=A;

		END IF;
	END PROCESS;
END A;
		
			
